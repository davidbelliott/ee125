library verilog;
use verilog.vl_types.all;
entity absolute_difference_vlg_vec_tst is
end absolute_difference_vlg_vec_tst;
