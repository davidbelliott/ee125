library verilog;
use verilog.vl_types.all;
entity log2_prob_vlg_vec_tst is
end log2_prob_vlg_vec_tst;
