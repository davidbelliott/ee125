-----------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
 
package user_types is
    type slv_array is array (natural range <>) of std_logic_vector;
end package;