library verilog;
use verilog.vl_types.all;
entity sync_counter_vlg_vec_tst is
end sync_counter_vlg_vec_tst;
