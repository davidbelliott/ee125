library verilog;
use verilog.vl_types.all;
entity leading_ones_sequential_vlg_vec_tst is
end leading_ones_sequential_vlg_vec_tst;
