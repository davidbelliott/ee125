library verilog;
use verilog.vl_types.all;
entity debouncer_demo_vlg_vec_tst is
end debouncer_demo_vlg_vec_tst;
